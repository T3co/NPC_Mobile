library ieee;
use ieee.std_logic_1164.all;
entity PWM_Controller is
port ( clk: in bit;  
       pOut : out STD_LOGIC);
end;
